module addRC (mem, cnt64_value, xor_en, slice);  //cnt_24 from full controller

    input [24:0] slice;
    input [5:0] cnt64_value;
    input xor_en;
    output reg [24:0] mem [63:0];  

    wire [7:0] cnt24_value; //badan input she

    assign cnt24_value = 8'd2;
    // reg [24:0] temp [63:0];
    
    reg [63:0] table_value;
    integer t_index;

    always @(posedge xor_en) begin  
        mem[cnt64_value] = slice;
        t_index = 63 - cnt64_value;
        mem[cnt64_value][12] = mem[cnt64_value][12] ^ table_value[t_index];          
    end

    always @(*) begin
        case(cnt24_value) 
            8'd00: table_value = 64'b0000000000000000000000000000000000000000000000000000000000000001;
            8'd01: table_value = 64'b0000000000000000000000000000000000000000000000001000000010000010;
            8'd02: table_value = 64'b1000000000000000000000000000000000000000000000001000000010001010;
            8'd03: table_value = 64'b1000000000000000000000000000000010000000000000001000000000000000;
            8'd04: table_value = 64'b0000000000000000000000000000000000000000000000001000000010001011;
            8'd05: table_value = 64'b0000000000000000000000000000000010000000000000000000000000000001;
            8'd06: table_value = 64'b1000000000000000000000000000000010000000000000001000000010000001;
            8'd07: table_value = 64'b1000000000000000000000000000000000000000000000001000000000001001;
            8'd08: table_value = 64'b0000000000000000000000000000000000000000000000000000000010001010;
            8'd09: table_value = 64'b0000000000000000000000000000000000000000000000000000000010001000;
            8'd10: table_value = 64'b0000000000000000000000000000000010000000000000001000000000001001;
            8'd11: table_value = 64'b0000000000000000000000000000000010000000000000000000000000001010;
            8'd12: table_value = 64'b0000000000000000000000000000000010000000000000001000000010001011;
            8'd13: table_value = 64'b1000000000000000000000000000000000000000000000000000000010001011;
            8'd14: table_value = 64'b1000000000000000000000000000000000000000000000001000000010001001;
            8'd15: table_value = 64'b1000000000000000000000000000000000000000000000001000000000000011;
            8'd16: table_value = 64'b1000000000000000000000000000000000000000000000001000000000000010;
            8'd17: table_value = 64'b1000000000000000000000000000000000000000000000000000000010000000;
            8'd18: table_value = 64'b0000000000000000000000000000000000000000000000001000000000001010;
            8'd19: table_value = 64'b1000000000000000000000000000000010000000000000000000000000001010;
            8'd20: table_value = 64'b1000000000000000000000000000000010000000000000001000000010000001;
            8'd21: table_value = 64'b1000000000000000000000000000000000000000000000001000000010000000;
            8'd22: table_value = 64'b0000000000000000000000000000000010000000000000000000000000000001;
            8'd23: table_value = 64'b1000000000000000000000000000000010000000000000001000000000001000;
        endcase
    end


endmodule