module datapath ();

endmodule


module controller ();

endmodule


module permutation_func ();

endmodule