module addRC (mem, cnt64_value, xor_en, slice, cnt24_value);  //cnt_24 from full controller

    input [24:0] slice;
    input [5:0] cnt64_value;
    input xor_en;
    output reg [24:0] mem [63:0];  

    input [4:0] cnt24_value; //badan input she

    // assign cnt24_value = 8'd0;
    // reg [24:0] temp [63:0];
    
    reg [63:0] table_value;
    integer t_index;

    always @(posedge xor_en) begin  
        mem[cnt64_value] = slice;
        t_index = 63 - cnt64_value;
        mem[cnt64_value][12] = mem[cnt64_value][12] ^ table_value[t_index];          
    end

    always @(*) begin
        case(cnt24_value) 
            5'd00: table_value = 64'b0000000000000000000000000000000000000000000000000000000000000001;
            5'd01: table_value = 64'b0000000000000000000000000000000000000000000000001000000010000010;
            5'd02: table_value = 64'b1000000000000000000000000000000000000000000000001000000010001010;
            5'd03: table_value = 64'b1000000000000000000000000000000010000000000000001000000000000000;
            5'd04: table_value = 64'b0000000000000000000000000000000000000000000000001000000010001011;
            5'd05: table_value = 64'b0000000000000000000000000000000010000000000000000000000000000001;
            5'd06: table_value = 64'b1000000000000000000000000000000010000000000000001000000010000001;
            5'd07: table_value = 64'b1000000000000000000000000000000000000000000000001000000000001001;
            5'd08: table_value = 64'b0000000000000000000000000000000000000000000000000000000010001010;
            5'd09: table_value = 64'b0000000000000000000000000000000000000000000000000000000010001000;
            5'd10: table_value = 64'b0000000000000000000000000000000010000000000000001000000000001001;
            5'd11: table_value = 64'b0000000000000000000000000000000010000000000000000000000000001010;
            5'd12: table_value = 64'b0000000000000000000000000000000010000000000000001000000010001011;
            5'd13: table_value = 64'b1000000000000000000000000000000000000000000000000000000010001011;
            5'd14: table_value = 64'b1000000000000000000000000000000000000000000000001000000010001001;
            5'd15: table_value = 64'b1000000000000000000000000000000000000000000000001000000000000011;
            5'd16: table_value = 64'b1000000000000000000000000000000000000000000000001000000000000010;
            5'd17: table_value = 64'b1000000000000000000000000000000000000000000000000000000010000000;
            5'd18: table_value = 64'b0000000000000000000000000000000000000000000000001000000000001010;
            5'd19: table_value = 64'b1000000000000000000000000000000010000000000000000000000000001010;
            5'd20: table_value = 64'b1000000000000000000000000000000010000000000000001000000010000001;
            5'd21: table_value = 64'b1000000000000000000000000000000000000000000000001000000010000000;
            5'd22: table_value = 64'b0000000000000000000000000000000010000000000000000000000000000001;
            5'd23: table_value = 64'b1000000000000000000000000000000010000000000000001000000000001000;
        endcase
    end


endmodule